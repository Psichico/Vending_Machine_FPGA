module vending_machine();


endmodule
